module str